module clockdivider (
	
);